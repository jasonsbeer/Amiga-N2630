----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:05:23 04/30/2022 
-- Design Name: 
-- Module Name:    U602 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity U602 is
    Port ( 
				A : IN  STD_LOGIC_VECTOR (31 downto 0);
				RnW : IN STD_LOGIC; --READ/WRITE SIGNAL FROM 680x0
				nAS : IN STD_LOGIC; --ADDRESS STROBE
				IORDY : IN STD_LOGIC; --IDE I/O READY
				INTRQ : IN STD_LOGIC; --IDE INTERUPT REQUEST
				MODE68K : IN STD_LOGIC; --ARE WE IN 68000 MODE?
				CPUCLK : IN STD_LOGIC; --25MHz CPU CLOCK
				nRESET : IN STD_LOGIC; --RESET SIGNAL
				IDEDIS : IN STD_LOGIC; --IDE DISABLE
				Z3DIS : IN STD_LOGIC; --ZORRO 3 RAM DISABLE
				nDS : IN STD_LOGIC; --68030 DATA STROBE
				FC : IN STD_LOGIC_VECTOR (2 DOWNTO 0); --68030 FUNCTION CODES
				SIZ : IN STD_LOGIC_VECTOR (1 DOWNTO 0); --68030 TRANSFER SIZE SIGNALS
				
				D : INOUT  STD_LOGIC_VECTOR (31 downto 24);
				
				nCS0 : OUT STD_LOGIC; --IDE CHIP SELECT 0
				nCS1 : OUT STD_LOGIC; --IDE CHIP SELECT 1
				DA : OUT STD_LOGIC_VECTOR (2 DOWNTO 0); --IDE ADDRESS LINES
				nDIOR : OUT STD_LOGIC; --IDE READ SIGNAL
				nDIOW : OUT STD_LOGIC; --IDE WRITE SIGNAL
				nDSACK0 : OUT STD_LOGIC; --68030 ASYNC PORT SIZE SIGNAL
				nDSACK1 : OUT STD_LOGIC; --68030 ASYNC PORT SIZE SIGNAL
				nDTACK : OUT STD_LOGIC; --68000 DATA SIGNAL
				nEM0UUBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, LOWER 64MB
				nEM0UMBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, LOWER 64MB
				nEM0LMBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, LOWER 64MB
				nEM0LLBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, LOWER 64MB
				nEM1UUBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, UPPER 64MB
				nEM1UMBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, UPPER 64MB
				nEM1LMBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, UPPER 64MB
				nEM1LLBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, UPPER 64MB
				EMA : OUT STD_LOGIC_VECTOR (12 DOWNTO 0); --ZORRO 3 MEMORY BUS
				BANK0 : OUT STD_LOGIC; --SDRAM BANK0
				BANK1 : OUT STD_LOGIC; --SDRAM BANK1
				nCAS0 : OUT STD_LOGIC;
				nRAS0 : OUT STD_LOGIC;
				nEM0WE : OUT STD_LOGIC;
				nEM0CS : OUT STD_LOGIC;
				EM0CLKE : OUT STD_LOGIC;				
				nCAS1 : OUT STD_LOGIC;
				nRAS1 : OUT STD_LOGIC;
				nEM1WE : OUT STD_LOGIC;
				nEM1CS : OUT STD_LOGIC;
				EM1CLKE : OUT STD_LOGIC;
				nSTERM : OUT STD_LOGIC
				
			);
end U602;

architecture Behavioral of U602 is

	SIGNAL IDE_SPACE : STD_LOGIC := '0'; --ARE WE IN THE IDE BASE ADDRESS SPACE?
	
	SIGNAL Z3RAM_BASE_ADDR : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL Z3RAM_CONFIGED : STD_LOGIC := '0'; --HAS ZORRO 3 RAM BEEN AUTOCONFIGed? ACTIVE HIGH
	SIGNAL Z3_AUTOCONFIG_SPACE :STD_LOGIC := '0'; --ARE WE IN THE ZORRO 3 AUTOCONFIG ADDRESS SPACE?
	
	SIGNAL DATAOUTAC : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => 'Z');
	SIGNAL DATAOUT : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => 'Z');
	
	SIGNAL MEMORY_SPACE : STD_LOGIC := '0'; --ARE WE IN THE ZORRO 3 MEMORY SPACE?
	SIGNAL LOW_MEMORY_SPACE : STD_LOGIC := '0'; --ACCESSING THE FIRST 64MB
	SIGNAL HIGH_MEMORY_SPACE : STD_LOGIC := '0'; --ADESSING THE SECOND 64MB
	
	--DEFINE THE SDRAM STATE MACHINE STATES
	TYPE SDRAM_STATE IS ( POWERUP, POWERUP_PRECHARGE, MODE_REGISTER, AUTO_REFRESH, AUTO_REFRESH_CYCLE, RUN_STATE, CAS_STATE, DATA_STATE );
	
	SIGNAL CURRENT_STATE : SDRAM_STATE;
	SIGNAL SDRAM_START_REFRESH_COUNT : STD_LOGIC := '0'; --WE NEED TO REFRESH TWICE UPON STARTUP	
	
	SIGNAL nUUBE : STD_LOGIC := '1'; --DYNAMIC BUS SIZE SIGNALS
	SIGNAL nUMBE : STD_LOGIC := '1';
	SIGNAL nLMBE : STD_LOGIC := '1';
	SIGNAL nLLBE : STD_LOGIC := '1';
	
	SIGNAL REFRESH_COUNTER : INTEGER RANGE 0 TO 255 := 0;
	SIGNAL COUNT : INTEGER RANGE 0 TO 2 := 0; --COUNTER FOR SDRAM STARTUP ACTIVITIES
	
	CONSTANT REFRESH_COUNTER_DEFAULT : INTEGER := 185;
	--AT 25MHZ, WE NEED TO REFRESH EVERY 195 CLOCK CYCLES
	--THIS CAUSES US TO REFRESH 8192 TIMES EVERY 64 MILLISECONDS
	--WE GO A LITTLE LESS THAN 195 IN CASE REFRESH HITS IN THE MIDDLE OF A RAM ACTION
	--THAT GIVES US SOME WIGGLE ROOM

begin

	---------------------
	-- DATA BUS OUTPUT --
	---------------------
	
	--WE ARE USING THE SAME DATA BITS IN SEVERAL PLACES.
	--THIS CREATES A SINGLE OUTPUT POINT, WHICH KEEPS VHDL HAPPY
	
	D(31 DOWNTO 24) <= 
			DATAOUTAC & "ZZZZ" WHEN Z3_AUTOCONFIG_SPACE = '1'
		ELSE 
			DATAOUT WHEN IDE_SPACE = '1'
		ELSE 
			"ZZZZZZZZ";

	----------------
	-- AUTOCONFIG --
	----------------
	
	--WE WILL AUTOCONFIG THE ZORRO 3 RAM (112MB) HERE
	--BECAUSE THIS IS IN THE ZORRO 3 SPACE, AUTOCONFIG IS DIFFERENT THAN THE ZORRO 2 AUTOCONFIG FOUND IN U601.
	--THE ZORRO 3 AUTCONFIG SPACE IS AT ADDRESS $FF00xxxx
	--WE ONLY AUTOCONFIG IF THE USER WANTS IT AND IT HAS NOT YET BEEN COMPLETED
	
	Z3_AUTOCONFIG_SPACE <= '1' WHEN A(31 DOWNTO 24) = x"FF" AND nAS = '0' AND Z3DIS = '1' AND Z3RAM_CONFIGED = '0' AND MODE68K = '0' ELSE '0';
	
	PROCESS (CPUCLK, nRESET) BEGIN
		
		IF nRESET = '0' THEN
			--COMPUTER HAS BEEN RESET
			Z3RAM_BASE_ADDR <= (OTHERS => '0');
			Z3RAM_CONFIGED <= '0';
		
		ELSIF RISING_EDGE(CPUCLK) THEN
			--START ZORRO 3 AUTOCONFIG
			IF Z3_AUTOCONFIG_SPACE = '1' THEN
				
				IF RnW = '1' THEN
					--READ REGISTERS
			
					CASE A(8 DOWNTO 2) IS
					
						--000
						--11111111000000000000000000000000
						WHEN "0000000" => DATAOUTAC <= "1010"; --zorro 3 card, link to system mem, not autoboot
						
						--100
						--11111111000000000000000100000000
						WHEN "1000000" => DATAOUTAC <= "0011"; --128mb		
						
						--004
						--11111111000000000000000000000100
						--WHEN "0000001" => D(31 DOWNTO 28) <= "1111"; --Product Number		
						
						--008
						--11111111000000000000000000001000
						--INVERTED
						WHEN "0000010" => DATAOUTAC <= "0000"; --Mem device, can't be shut up
						
						--108
						--11111111000000000000000100001000
						--INVERTED
						WHEN "1000010" => DATAOUTAC <= "1110"; --Automatically sized by the OS						
					
						WHEN OTHERS => DATAOUTAC <= "1111";
					
					END CASE;
					
				ELSE
					--WRITE REGISTER
					
					--44
					--11111111000000000000000001000100.
					--THIS IS THE BASE ADDRESS OF THE Z3 RAM
					IF A(8 DOWNTO 2) = "0010001" AND nDS = '0' THEN				
						
						Z3RAM_BASE_ADDR <= D(31 DOWNTO 27);
						Z3RAM_CONFIGED <= '1';
						
					END IF;
					
				END IF;
			
			END IF;
		END IF;
	END PROCESS;


	------------------------------------------------------
	-- GAYLE COMPATABLE HARD DRIVE CONTROLLER INTERFACE --
	------------------------------------------------------

	--WE ARE GOING TO USE THE AMIGA OS GAYLE IDE INTERFACE
	--UNFORTUNATELY, THIS MEANS VERY LIMITED PERFORMANCE CAPABILITY, ONLY SUPPORTING PIO 0 WITH UP TO 2 DRIVES.
	--BUT IT IS SIMPLE TO IMPLEMENT AND READY OUT OF THE BOX WITH KS 35.300.
	--COMPATABILITY CAN BE ADDED TO EARLIER KICKSTARTS BY ADDING THE APPROPRIATE SCSI.DEVICE TO ROM
	--IN THE FUTURE, I WOULD LIKE TO REPLACE THIS WITH A MORE ROBUST MULTIDRIVE IDE INTERFACE
	
	--GAYLE IS ONLY CONNECTED TO A23..12, SO WE ARE IMITATING THAT HERE

	--TO TRICK AMIGA OS INTO THINKING WE HAVE A GAYLE ADDRESS DECODER, WE NEED TO RESPOND TO GAYLE SPECIFIC REGISTERS
	--SEE THE GAYLE SPECIFICATIONS FOR MORE DETAILS.
	--WE DISABLE THE IDE PORT BY SIMPLY IGNORING THE GAYLE CONFIGURATION REGISTERS, WHICH TELLS AMIGA OS THERE IS NO GAYLE HERE.
	
	--IN THE EVENT THE IDE DEVICE IS ASSERTING AN INTERRUPT REQUEST, WE PASS THAT TO ANYONE INTERESTED WITH THE REGISTER AT $DA8000.
	--BIT 7 IS SET HIGH TO INDICATE THE IRQ. THE OTHER BITS ARE ALL FOR THE PCMCIA, SETTING BIT 0 HIGH DISABLES IT.
	--THE INTERUPT REQUEST IS ACKNOWLEDGED WITH THE REGISTER AT $DA9000. THERE IS NOT A HARDWARE INTERUPT ACK, SO JUST FYI.	
	
	PROCESS (CPUCLK) BEGIN
		IF (RISING_EDGE (CPUCLK)) THEN
		
			IF (RnW = '1' AND nAS = '0' AND IDEDIS = '1') THEN
			
				CASE A(23 DOWNTO 12) IS
					WHEN x"DE1" => DATAOUT <= x"DF"; --GAYLE_ID is at $DE1000. Return $DF.
					WHEN x"DAA" => DATAOUT <= x"80"; --INTENA (enable ide interupts) AT $DAA000, Return $80.
					WHEN x"DA8" => DATAOUT <= INTRQ & "0000001"; --IDE Device Interrupt Request on data bit 7 at $DA8000.
					WHEN OTHERS => DATAOUT <= (OTHERS => 'Z');
				END CASE;
				
			END IF;
			
		END IF;
	END PROCESS;
	
	--GAYLE SPECS TELL US WHEN THE IDE CHIP SELECT LINES ARE ACTIVE
	
	nCS0 <= '0' 
		WHEN 
			(A(14 DOWNTO 12) = "000" OR A(14 DOWNTO 12) = "010") AND nAS = '0' --$0DA0000 TO $0DA0FFF OR $0DA2000 TO $0DA2FFF
		ELSE 
			'1';
			
	nCS1 <= '0' 
		WHEN 
			(A(14 DOWNTO 12) = "001" OR A(14 DOWNTO 12) = "011") AND nAS = '0' --$0DA1000 TO $0DA1FFF OR $0DA3000 TO $0DA3FFF
		ELSE 
			'1';
			
	--GAYLE EXPECTS IDE DA2..0 TO BE CONNECTED TO A4..2
	
	DA(0) <= A(2);
	DA(1) <= A(3);
	DA(2) <= A(4);
	
	--ARE WE IN THE ASSIGNED ADDRESS SPACE FOR THE IDE CONTROLLER?
	--GAYLE IDE ADDRESS SPACE IS $0DA0000 - $0DA3FFF. THE ADDRESS SPACE IS HARD CODED.
	--SPACE $0DA4000 - $0DA4FFF IS IDE RESERVED. GUESSING IT WAS NEVER IMPLEMENTED? MAYBE FOR A SECOND PORT?
	IDE_SPACE <= '1' WHEN (A(23 DOWNTO 12) >= x"DA0" AND A(23 DOWNTO 12) <= x"DA3") AND nAS = '0' ELSE '0';
	
	--HERE IS THE CONTROLLER INTERFACE
	PROCESS (CPUCLK, nRESET) BEGIN
	
		IF (nRESET = '0') THEN
			--AMIGA HAS RESET, START OVER
			nDIOR <= '1';
			nDIOW <= '1';
			nDSACK0 <= 'Z';
			nDSACK1 <= 'Z';
			nDTACK <= 'Z';
		
		ELSIF (RISING_EDGE(CPUCLK)) THEN
		
			IF (IDE_SPACE = '1') THEN			
				--WE ARE IN THE IDE ADDRESS SPACE 
				
				 IF (nAS = '0') THEN 
					--ADDRESS STROBE IS ASSERTED
				
					IF (RnW = '1') THEN
						--THIS IS A READ
						nDIOR <= '0';
						nDIOW <= '1';
					ELSE
						--THIS IS A WRITE
						nDIOR <= '1';
						nDIOW <= '0';
					END IF;
						
					IF (IORDY = '1') THEN
					
						--THE DEVICE IS READY TO TRANSMIT OR RECEIVE DATA, SIGNAL 16 BIT PORT TO 68030
						--DTACK WHEN IN 68K MODE
						IF (MODE68K = '0') THEN
							nDSACK0 <= '1';
							nDSACK1 <= '0';
						ELSE
							nDTACK <= '0';
						END IF;
						
					END IF;
					
				ELSE
				
					--ADDRESS STROBE NOT ASSERTED
					IF (MODE68K = '0') THEN
						nDSACK0 <= '1';
						nDSACK1 <= '1';
					ELSE
						nDTACK <= '1';
					END IF;
					
				END IF;	
			
			ELSE
			
				--SET IN A "NOP" STATE
				nDIOR <= '1';
				nDIOW <= '1';
				
				--HI Z DSACK/DTACK SO WE DON'T INTERFERE WITH OTHER STUFF ON THE BUS
				IF (MODE68K = '0') THEN
					nDSACK0 <= 'Z';
					nDSACK1 <= 'Z';
				ELSE
					nDTACK <= 'Z';
				END IF;
					
			END IF;
		
		END IF;
	
	END PROCESS;

	------------------------------
	-- ZORRO 3 MEMORY CONTROLER --
	------------------------------
	
	--ARE WE ACCESSING THE Z3 MEMORY?
	MEMORY_SPACE <= '1' WHEN 
			A(31 DOWNTO 27) = Z3RAM_BASE_ADDR AND nAS = '0' AND Z3RAM_CONFIGED = '1' AND FC(2 DOWNTO 0) = "111" 
		ELSE 
			'0';

	--DETERMINE WHAT SPACE IN THE MEMORY WE ARE ACCESSING
	--THIS DETERMINES WHICH PAIR OF SDRAMS WE ARE ACCESSING
	LOW_MEMORY_SPACE <= '1' WHEN A(26) = '0' AND MEMORY_SPACE = '1' ELSE '0';
	HIGH_MEMORY_SPACE <= '1' WHEN A(26) = '1' AND MEMORY_SPACE = '1' ELSE '0';
	
	--SET THE DYNAMIC BUS SIZING
	nEM0UUBE <= nUUBE;
	nEM0UMBE <= nUMBE;
	nEM0LMBE <= nLMBE;
	nEM0LLBE <= nLLBE;
	
	nEM1UUBE <= nUUBE;
	nEM1UMBE <= nUMBE;
	nEM1LMBE <= nLMBE;
	nEM1LLBE <= nLLBE;
	
	-------------------------------------
	-- SDRAM FALLING CLOCK EDGE ACTIONS --
	-------------------------------------
	
	PROCESS ( CPUCLK ) BEGIN
		
		IF ( FALLING_EDGE (CPUCLK) ) THEN

			IF (MEMORY_SPACE = '1') THEN		

				--ENABLE THE VARIOUS BYTES ON THE SDRAM DEPENDING ON WHAT THE ACCESSING DEVICE IS ASKING FOR. U603
				--DISCUSSION OF PORT SIZE AND BYTE SIZING IS ALL IN SECTION 12 OF THE 68030 USER MANUAL.
				
				--UPPER UPPER BYTE ENABLE (D31..24)
				IF 
				   (( RnW = '1' ) OR
					(A(1 downto 0) = "00" AND nDS = '0'))
				THEN			
					nUUBE <= '0'; 
				ELSE 
					nUUBE <= '1';
				END IF;

				--UPPER MIDDLE BYTE (D23..16)
				IF 
					(( RnW = '1' ) OR
					(A(1 downto 0) = "01" AND nDS = '0') OR
					(A(1) = '0' AND SIZ(0) = '0'  AND nDS = '0') OR
					(A(1) = '0' AND SIZ(1) = '1'  AND nDS = '0')) 
				THEN
					nUMBE <= '0';
				ELSE
					nUMBE <= '1';
				END IF;

				--LOWER MIDDLE BYTE (D15..8)
				IF 
				   (( RnW = '1' ) OR
					(A(1 downto 0) = "10" AND nDS = '0') OR
					(A(1) = '0' AND SIZ(0) = '0' AND SIZ(1) = '0'  AND nDS = '0') OR
					(A(1) = '0' AND SIZ(0) = '1' AND SIZ(1) = '1'  AND nDS = '0') OR
					(A(0) = '1' AND A(1) = '0' AND SIZ(0) = '0'  AND nDS = '0'))
				THEN
					nLMBE <= '0';
				ELSE
					nLMBE <= '1';
				END IF;

				--LOWER LOWER BYTE (D7..0)
				IF 
				   (( RnW = '1' ) OR
					(A(1 downto 0) = "11" AND nDS = '0' ) OR
					(A(0) = '1' AND SIZ(0) = '1' AND SIZ(1) = '1' AND nDS = '0') OR
					(SIZ(0) = '0' AND SIZ(1) = '0' AND nDS = '0') OR
					(A(1) = '1' AND SIZ(1) ='1' AND nDS = '0'))
				THEN
					nLLBE <= '0';
				ELSE
					nLLBE <= '1';
				END IF;	

			ELSE 
				--DEACTIVATE ALL THE RAM BYTE MASKS

				nUUBE <= '1';
				nUMBE <= '1';
				nLMBE <= '1';
				nLLBE <= '1';

			END IF;	
		END IF;
	END PROCESS;
	
	
	-------------------------------------
	-- SDRAM RISING CLOCK EDGE ACTIONS --
	-------------------------------------
	
	PROCESS ( CPUCLK, nRESET ) BEGIN
	
		IF (nRESET = '0') THEN 
				--THE AMIGA HAS BEEN RESET
				CURRENT_STATE <= POWERUP;
				
				nCAS0 <= '1';
				nRAS0 <= '1';
				nEM0WE <= '1';
				nEM0CS <= '1';
				EM0CLKE <= '0';
				
				nCAS1 <= '1';
				nRAS1 <= '1';
				nEM1WE <= '1';
				nEM1CS <= '1';
				EM1CLKE <= '0';
				
				COUNT <= 0;
				SDRAM_START_REFRESH_COUNT <= '0';
				nSTERM <= 'Z';
				
		ELSIF ( RISING_EDGE (CPUCLK) ) THEN
			
			--SDRAM is pretty fast. Most operations will complete in less than one 25MHz clock cycle. Only AUTOREFRESH and 
			--successive BANK ACTIVE commands take more than one clock cycle. Both are 60ns.
			
			--REFRESH
			IF (REFRESH_COUNTER >= REFRESH_COUNTER_DEFAULT) THEN
				--TIME TO REFRESH THE SDRAM
				IF (MEMORY_SPACE = '0') THEN
					--IF THIS IS NOT A MEMORY CYCLE, PROCEED DIRECTLY TO REFRESH
					--IF WE ARE IN THE MIDDLE OF MEMORY ACCESS, WE NEED TO WAIT UNTIL THAT IS OVER
					CURRENT_STATE <= AUTO_REFRESH;
				END IF;
			ELSE
				--INCREMENT THE REFRESH COUNTER
				REFRESH_COUNTER <= REFRESH_COUNTER + 1;
			END IF;
		
			--PROCEED WITH SDRAM STATE MACHINE
			--THE FIRST STATES ARE TO INITIALIZE THE SDRAM, WHICH WE ALWAYS DO
			--THE LATER STATES ARE TO UTILIZE THE SDRAM, WHICH ONLY HAPPENS IF MEMORY_SPACE = 1
			--THIS MEANS THE ADDRESS STROBE IS ASSERTED, WE ARE IN THE ZORRO 3 ADDRESS SPACE, AND THE RAM IS AUTOCONFIGured
			CASE CURRENT_STATE IS
			
				WHEN POWERUP =>
					--First power up or warm reset
					--200 microsecond is needed to stabilize. We are going to rely on the 
					--the system reset to give us the needed time, although it might be inadequate.
					
					nCAS0 <= '1';
					nRAS0 <= '1';
					nEM0WE <= '1';
					nEM0CS <= '1';
					EM0CLKE <= '0';
					
					nCAS1 <= '1';
					nRAS1 <= '1';
					nEM1WE <= '1';
					nEM1CS <= '1';
					EM1CLKE <= '0';
					
					CURRENT_STATE <= POWERUP_PRECHARGE;
					
				WHEN POWERUP_PRECHARGE =>
					--ALL BANKS TO BE PRECHARGED
					EMA <= (OTHERS => '0');
					EMA(10) <= '1'; --PRECHARGE ALL	
					
					nCAS0 <= '1';
					nRAS0 <= '0';
					nEM0WE <= '0';
					nEM0CS <= '0';
					nEM0CLKE <= '1';
					
					nCAS1 <= '1';
					nRAS1 <= '0';
					nEM1WE <= '0';
					nEM1CS <= '0';
					nEM1CLKE <= '1';
					
					CURRENT_STATE <= MODE_REGISTER;
				
				WHEN MODE_REGISTER =>
					--TWO CLOCK CYCLES ARE NEEDED FOR THE REGISTER TO, WELL, REGISTER
					EMA <= "0001000100000"; --PROGRAM THE SDRAM...NO READ OR WRITE BURST, CAS LATENCY=2,
					
					nCAS0 <= '0';
					nRAS0 <= '0';
					nEM0WE <= '0';
					nEM0CS <= '0';
					
					nCAS1 <= '0';
					nRAS1 <= '0';
					nEM1WE <= '0';
					nEM1CS <= '0';
					
					IF (COUNT = 1) THEN
						--NOW NEED TO REFRESH TWICE
						CURRENT_STATE <= AUTO_REFRESH;
					END IF;
					
					COUNT <= COUNT + 1;
					
				WHEN AUTO_REFRESH =>
					--REFRESH the SDRAM
					--MUST BE FOLLOWED BY NOPs UNTIL REFRESH COMPLETE
					--Refresh time is 60ns. Each 25MHz clock period is 40ns.
					--If we wait two clock cycles, this will allow time for refresh.
					
					nCAS0 <= '0';
					nRAS0 <= '0';
					nEM0WE <= '1';
					nEM0CS <= '0';
					
					nCAS1 <= '0';
					nRAS1 <= '0';
					nEM1WE <= '1';
					nEM1CS <= '0';					
					
					COUNT <= 0;
					
					CURRENT_STATE <= AUTO_REFRESH_CYCLE;				
					
				WHEN AUTO_REFRESH_CYCLE =>
					--NOPs WHILE THE SDRAM IS REFRESHING
					
					nCAS0 <= '1';
					nRAS0 <= '1';
					nEM0WE <= '1';
					nEM0CS <= '1';
					
					nCAS1 <= '1';
					nRAS1 <= '1';
					nEM1WE <= '1';
					nEM1CS <= '1';	
					
					IF (COUNT = 1) THEN --TWO CLOCK CYCLES HAVE PASSED. WE CAN PROCEED.
						--DO WE NEED TO REFRESH AGAIN (STARTUP)?
						IF (SDRAM_START_REFRESH_COUNT = '0') THEN							
							CURRENT_STATE <= AUTO_REFRESH;
							SDRAM_START_REFRESH_COUNT <= '1';
						ELSE
							--DESELECT ALL SDRAMs
							nEM0CS <= '1';
							nEM1CS <= '1';	
							
							--WE SHOULD BE READY TO GO!
							CURRENT_STATE <= RUN_STATE;
							REFRESH_COUNTER <= 0;
						END IF;
					END IF;		

					COUNT <= COUNT + 1;						
				
				WHEN RUN_STATE =>
					--CLOCK EDGE 0
					
					IF (MEMORY_SPACE = '1') THEN 
						--WE ARE IN THE Z3 MEMORY SPACE WITH THE ADDRESS STROBE ASSERTED.
						--SEND THE BANK ACTIVATE COMMAND W/RAS
						
						--SELECT THE CORRECT SET OF SDRAMs BASED ON ADDRESS
						IF (LOW_MEMORY_SPACE = '1') THEN nEM0CS <= '0'; ELSE nEM0CS <= '1'; END IF;
						IF (HIGH_MEMORY_SPACE = '1') THEN nEM1CS <= '0'; ELSE nEM1CS <= '1'; END IF;
						
						EMA(12 downto 0) <= A(14 downto 2);
						BANK0 <= A(15);
						BANK1 <= A(16);
						
						--HERE, I'M SENDING THE COMMANDS TO ALL SDRAMs, BUT ONLY THE SELECTED PAIR SHOULD RESPOND
						nCAS0 <= '1';
						nRAS0 <= '0';
						nEM0WE <= '1';
						
						nCAS1 <= '1';
						nRAS1 <= '0';
						nEM1WE <= '1';
						
						nSTERM <= '1'; --WE ARE USING THE BUS RIGHT NOW, SO NEGATE STERM IN PREPARTATION FOR USE
						
						CURRENT_STATE <= CAS_STATE;
						COUNT <= 0;
					END IF;
					
				WHEN CAS_STATE =>
					--CLOCK EDGE 1
					--READ OR WRITE WITH AUTOPRECHARGE
					
					EMA(8 downto 0) <= A(25 downto 17);
					EMA(9) <= '0';
					EMA(10) <= '1'; --AUTO PRECHARGE
					
					nCAS0 <= '0';
					nRAS0 <= '1';
					nEM0WE <= RnW;
					
					nCAS1 <= '0';
					nRAS1 <= '1';
					nEM1WE <= RnW;

					--IF THIS IS A WRITE ACTION, WE CAN IMMEDIATELY PROCEED TO THE ACTION
					--IF THIS IS A READ ACTION, THE CAS LATENCY IS 2 CLOCK CYCLES, SO WE NEED TO WAIT ONE MORE CLOCK BEFORE READING
					--DURING DMA, THE REQUESTING DEVICE'S RW SIGNAL IS LOCKED TO OUR RW SIGNAL

					IF ((RnW = '0') OR (RnW = '1' AND COUNT >= 1)) THEN
					
						nSTERM <= '0';
						
						CURRENT_STATE <= DATA_STATE;
					
					END IF;						
					
					COUNT <= COUNT + 1;
					
				WHEN DATA_STATE =>
					--RISING CLOCK EDGE 2
					--THIS IS THE CLOCK EDGE WE EXPECT THE DATA TO BE WRITTEN TO OR READ FROM THE SDRAM
					--WE NEED TO WAIT 30ns BEFORE ISSUING ANOTHER BANK ACTIVATE COMMAND. NO PROBLEM, SINCE ONE CLOCK CYCLE IS 40ns.
					
					IF (MEMORY_SPACE = '0') THEN --THE ADDRESS STROBE HAS NEGATED INDICATING THE END OF THE MEMORY ACCESS
						
						--TRISTATE SO WE DON'T INTERFERE WITH OTHER DEVICES ON THE BUSES
						nSTERM <= 'Z';
						
						CURRENT_STATE <= RUN_STATE;
						
						--SET NOP
						nCAS0 <= '1';
						nRAS0 <= '1';
						nEM0WE <= '1';
						nEM0CS <= '1';
						
						nCAS1 <= '1';
						nRAS1 <= '1';
						nEM1WE <= '1';
						nEM1CS <= '1';
						
					END IF;					
				
			END CASE;
				
		END IF;
	END PROCESS;

end Behavioral;

