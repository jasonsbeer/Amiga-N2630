--This work is shared under the Attribution-NonCommercial-ShareAlike 4.0 International (CC BY-NC-SA 4.0) License
--https://creativecommons.org/licenses/by-nc-sa/4.0/legalcode
	
--You are free to:
--Share - copy and redistribute the material in any medium or format
--Adapt - remix, transform, and build upon the material

--Under the following terms:

--Attribution - You must give appropriate credit, provide a link to the license, and indicate if changes were made. 
--You may do so in any reasonable manner, but not in any way that suggests the licensor endorses you or your use.

--NonCommercial - You may not use the material for commercial purposes.

--ShareAlike - If you remix, transform, or build upon the material, you must distribute your contributions under the 
--same license as the original.

--No additional restrictions - You may not apply legal terms or technological measures that legally restrict others 
--from doing anything the license permits.

----------------------------------------------------------------------------------
-- Company: 
-- Engineer:       JASON NEUS
-- 
-- Create Date:    09:42:54 02/13/2022 
-- Design Name:    N2630 U602 CPLD
-- Module Name:    U600 - Behavioral 
-- Project Name:   N2630
-- Target Devices: XC95144 144 PIN
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 1.0 - Original Release
-- Additional Comments: EQUATIONS FOR THE N2630 PROJECT BY JASON NEUS.
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity U602 is
    Port ( 
				A : IN  STD_LOGIC_VECTOR (31 downto 0);
				RnW : IN STD_LOGIC; --READ/WRITE SIGNAL FROM 680x0
				nAS : IN STD_LOGIC; --ADDRESS STROBE
				IORDY : IN STD_LOGIC; --IDE I/O READY
				INTRQ : IN STD_LOGIC; --IDE INTERUPT REQUEST
				MODE68K : IN STD_LOGIC; --ARE WE IN 68000 MODE?
				CPUCLK : IN STD_LOGIC; --25MHz CPU CLOCK
				nRESET : IN STD_LOGIC; --SYSTEM RESET SIGNAL VALID IN 68000 AND 68030 MODE
				nGRESET : IN STD_LOGIC; --68030 ONLY RESET SIGNAL
				nIDEDIS : IN STD_LOGIC; --IDE DISABLE
				nZ3DIS : IN STD_LOGIC; --ZORRO 3 RAM DISABLE
				nDS : IN STD_LOGIC; --68030 DATA STROBE
				FC : IN STD_LOGIC_VECTOR (2 DOWNTO 0); --68030 FUNCTION CODES
				SIZ : IN STD_LOGIC_VECTOR (1 DOWNTO 0); --68030 TRANSFER SIZE SIGNALS
				nBGACK : IN STD_LOGIC; --680x0 BUS GRANT ACK
	    			--SPEED : IN STD_LOGIC_VECTOR (1 DOWNTO 0); --USER SELECTED SDRAM REFRESH SPEED
				
				D : INOUT  STD_LOGIC_VECTOR (31 downto 24);
				EXTSEL : INOUT STD_LOGIC; --SIGNALS THE OTHER LOGIC THAT WE ARE RESPONDING TO THE RAM ADDRESS SPACE
				
				nCS0 : OUT STD_LOGIC; --IDE CHIP SELECT 0
				nCS1 : OUT STD_LOGIC; --IDE CHIP SELECT 1
				DA : OUT STD_LOGIC_VECTOR (2 DOWNTO 0); --IDE ADDRESS LINES
				nDIOR : OUT STD_LOGIC; --IDE READ SIGNAL
				nDIOW : OUT STD_LOGIC; --IDE WRITE SIGNAL
				--nDSACK0 : OUT STD_LOGIC; --68030 ASYNC PORT SIZE SIGNAL
				nDSACK1 : OUT STD_LOGIC; --68030 ASYNC PORT SIZE SIGNAL
				nDTACK : OUT STD_LOGIC; --68000 DATA SIGNAL
				nEM0UUBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, LOWER 64MB
				nEM0UMBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, LOWER 64MB
				nEM0LMBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, LOWER 64MB
				nEM0LLBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, LOWER 64MB
				nEM1UUBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, UPPER 64MB
				nEM1UMBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, UPPER 64MB
				nEM1LMBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, UPPER 64MB
				nEM1LLBE : OUT STD_LOGIC; --68030 DYNAMIC BUS SIZING OUTPUT, UPPER 64MB
				EMA : OUT STD_LOGIC_VECTOR (12 DOWNTO 0); --ZORRO 3 MEMORY BUS
				BANK0 : OUT STD_LOGIC; --SDRAM BANK0
				BANK1 : OUT STD_LOGIC; --SDRAM BANK1
				nCAS0 : OUT STD_LOGIC; --CAS LOW BANK
				nRAS0 : OUT STD_LOGIC; --RAS LOW BANK
				nEM0WE : OUT STD_LOGIC; --WRITE ENABLE LOW BANK
				nEM0CS : OUT STD_LOGIC; --CHIP SELECT LOW BANK
				EM0CLKE : OUT STD_LOGIC; --CLOCK ENABLE LOW BANK
				nCAS1 : OUT STD_LOGIC; --CAS HIGH BANK
				nRAS1 : OUT STD_LOGIC; --RAS HIGH BANK
				nEM1WE : OUT STD_LOGIC; --WRITE ENABLE HIGH BANK
				nEM1CS : OUT STD_LOGIC; --CHIP SELECT HIGH BANK
				EM1CLKE : OUT STD_LOGIC; --CLOCK ENABLE HIGH BANK
				nSTERM : OUT STD_LOGIC --68030 SYNCRONOUS TERMINATION SIGNAL
				
			);
end U602;

architecture Behavioral of U602 is

	SIGNAL IDE_SPACE : STD_LOGIC := '0'; --ARE WE IN THE IDE BASE ADDRESS SPACE?
	
	SIGNAL Z3RAM_BASE_ADDR : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL Z3RAM_CONFIGED : STD_LOGIC := '0'; --HAS ZORRO 3 RAM BEEN AUTOCONFIGed? ACTIVE HIGH
	SIGNAL Z3_AUTOCONFIG_SPACE :STD_LOGIC := '0'; --ARE WE IN THE ZORRO 3 AUTOCONFIG ADDRESS SPACE?
	
	SIGNAL DATAOUTAC : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => 'Z');
	SIGNAL DATAOUT : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => 'Z');
	
	SIGNAL MEMORY_SPACE : STD_LOGIC := '0'; --ARE WE IN THE ZORRO 3 MEMORY SPACE?
	SIGNAL LOW_MEMORY_SPACE : STD_LOGIC := '0'; --ACCESSING THE FIRST 64MB
	SIGNAL HIGH_MEMORY_SPACE : STD_LOGIC := '0'; --ADESSING THE SECOND 64MB
	
	--DEFINE THE SDRAM STATE MACHINE STATES
	TYPE SDRAM_STATE IS ( POWERUP, POWERUP_PRECHARGE, MODE_REGISTER, AUTO_REFRESH, AUTO_REFRESH_CYCLE, RUN_STATE, CAS_STATE, DATA_STATE );
	
	SIGNAL CURRENT_STATE : SDRAM_STATE;
	SIGNAL SDRAM_START_REFRESH_COUNT : STD_LOGIC := '0'; --WE NEED TO REFRESH TWICE UPON STARTUP	
	
	SIGNAL nUUBE : STD_LOGIC := '1'; --DYNAMIC BUS SIZE SIGNALS
	SIGNAL nUMBE : STD_LOGIC := '1';
	SIGNAL nLMBE : STD_LOGIC := '1';
	SIGNAL nLLBE : STD_LOGIC := '1';
	
	SIGNAL REFRESH_COUNTER : INTEGER RANGE 0 TO 255 := 0;
	SIGNAL COUNT : INTEGER RANGE 0 TO 3 := 0; --COUNTER FOR SDRAM STARTUP ACTIVITIES
	
	--CONSTANT REFRESH_COUNTER_25 : INTEGER := 185;
	--CONSTANT REFRESH_COUNTER_33 : INTEGER := 244;
	--CONSTANT REFRESH_COUNTER_40 : INTEGER := 296;
	--CONSTANT REFRESH_COUNTER_50 : INTEGER := 370;

	CONSTANT REFRESH_COUNTER_DEFAULT : INTEGER := 185; --25MHz
	--AT 25MHZ, WE NEED TO REFRESH EVERY 195 CLOCK CYCLES
	--THIS CAUSES US TO REFRESH 8192 TIMES EVERY 64 MILLISECONDS
	--WE GO A LITTLE LESS THAN 195 IN CASE REFRESH HITS IN THE MIDDLE OF A RAM ACTION
	--THAT GIVES US SOME WIGGLE ROOM

begin
	-------------------------
	-- AUTOREFRESH COUNTER --
	-------------------------
	
	--SET THE REFRESH COUNTER TO THE NUMBER SPECIFIED BY THE USER VIA JUMPERS	
	--CASE SPEED (1 DOWNTO 0) IS
		
		--WHEN "00" => CONSTANT REFRESH_COUNTER_DEFAULT <= REFRESH_COUNTER_50; --50MHz
		--WHEN "01" => CONSTANT REFRESH_COUNTER_DEFAULT <= REFRESH_COUNTER_40; --40MHz
		--WHEN "10" => CONSTANT REFRESH_COUNTER_DEFAULT <= REFRESH_COUNTER_33; --33MHz
		--WHEN "11" => CONSTANT REFRESH_COUNTER_DEFAULT <= REFRESH_COUNTER_25; --25MHz
			
	--END CASE;

	---------------------
	-- DATA BUS OUTPUT --
	---------------------
	
	--WE ARE USING THE SAME DATA BITS IN SEVERAL PLACES.
	--THIS CREATES A SINGLE OUTPUT POINT, WHICH KEEPS EVERYTHING HAPPY
	
	D(31 DOWNTO 24) <= 
			DATAOUTAC & "ZZZZ" WHEN Z3_AUTOCONFIG_SPACE = '1'
		ELSE 
			DATAOUT;

	----------------
	-- AUTOCONFIG --
	----------------
	
	--WE AUTOCONFIG THE ZORRO 3 RAM (UP TO 256MB) HERE
	--BECAUSE THIS IS IN THE ZORRO 3 SPACE, AUTOCONFIG IS DIFFERENT THAN THE ZORRO 2 AUTOCONFIG FOUND IN U601.
	--THE ZORRO 3 AUTCONFIG SPACE IS AT ADDRESS $FF00xxxx
	--WE ONLY AUTOCONFIG IF THE 68030 IS NOT IN RESET, THE USER WANTS IT, AND IT HAS NOT YET BEEN COMPLETED
	--WE AUTOCONFIG HERE BECAUSE THE EXTRA RAM IS TECHNICALLY OPTIONAL.
	
	Z3_AUTOCONFIG_SPACE <= '1' WHEN A(31 DOWNTO 24) = x"FF" AND nAS = '0' AND nZ3DIS = '1' AND Z3RAM_CONFIGED = '0' ELSE '0';
	
	PROCESS (CPUCLK, nGRESET) BEGIN
		
		IF nGRESET = '0' THEN
			--68030 HAS BEEN RESET
			Z3RAM_CONFIGED <= '0';
		
		ELSIF RISING_EDGE(CPUCLK) THEN
			--START ZORRO 3 AUTOCONFIG
			IF Z3_AUTOCONFIG_SPACE = '1' THEN
				
				IF RnW = '1' THEN
					--READ REGISTERS
			
					CASE A(8 DOWNTO 2) IS
					
						--000
						--11111111000000000000000000000000
						WHEN "0000000" => DATAOUTAC <= "1010"; --zorro 3 card, link to system mem, not autoboot
						
						--100
						--11111111000000000000000100000000
						WHEN "1000000" => DATAOUTAC <= "0011"; --128mb		
						
						--004
						--11111111000000000000000000000100
						--WHEN "0000001" => D(31 DOWNTO 28) <= "1111"; --Product Number		
						
						--008
						--11111111000000000000000000001000
						--INVERTED
						WHEN "0000010" => DATAOUTAC <= "0000"; --Mem device, can't be shut up
						
						--108
						--11111111000000000000000100001000
						--INVERTED
						WHEN "1000010" => DATAOUTAC <= "1110"; --Automatically sized by the OS						
					
						WHEN OTHERS => DATAOUTAC <= "1111";
					
					END CASE;
					
				ELSE
					--WRITE REGISTER
					
					--44
					--11111111000000000000000001000100.
					--THIS IS THE BASE ADDRESS OF THE Z3 RAM
					IF A(8 DOWNTO 2) = "0010001" AND nDS = '0' THEN				
						
						Z3RAM_BASE_ADDR <= D(31 DOWNTO 27);
						Z3RAM_CONFIGED <= '1';
						
					END IF;
					
				END IF;
			
			END IF;
		END IF;
	END PROCESS;


	------------------------------------------------------
	-- GAYLE COMPATABLE HARD DRIVE CONTROLLER INTERFACE --
	------------------------------------------------------

	--WE ARE GOING TO USE THE AMIGA OS GAYLE IDE INTERFACE
	--UNFORTUNATELY, THIS MEANS ONLY SUPPORTING PIO WITH UP TO 2 DRIVES.
	--BUT IT IS SIMPLE TO IMPLEMENT AND READY OUT OF THE BOX WITH KS => 35.300.
	--COMPATABILITY CAN BE ADDED TO EARLIER KICKSTARTS BY ADDING THE APPROPRIATE SCSI.DEVICE TO ROM
	--IN THE FUTURE, I WOULD LIKE TO REPLACE THIS WITH A MORE ROBUST MULTIPORT IDE INTERFACE PREFERABLY WITH DMA.
			
	--PERFORMACE SHOULD BE RESPECTABLE WITH THE 68030, BUT ANEMIC IN 68000 MODE.
	
	--GAYLE IS ONLY CONNECTED TO A23..12, SO WE ARE IMITATING THAT HERE

	--TO TRICK AMIGA OS INTO THINKING WE HAVE A GAYLE ADDRESS DECODER, WE NEED TO RESPOND TO GAYLE SPECIFIC REGISTERS
	--SEE THE GAYLE SPECIFICATIONS FOR MORE DETAILS.
	--WE DISABLE THE IDE PORT BY SIMPLY IGNORING THE GAYLE CONFIGURATION REGISTERS, WHICH TELLS AMIGA OS THERE IS NO GAYLE HERE.
	
	--IN THE EVENT THE IDE DEVICE IS ASSERTING AN INTERRUPT REQUEST, WE PASS THAT TO ANYONE INTERESTED WITH THE REGISTER AT $DA8000.
	--BIT 7 IS SET HIGH TO INDICATE THE IRQ. THE OTHER BITS ARE ALL FOR THE PCMCIA, SETTING BIT 0 HIGH DISABLES IT.
	--THE INTERUPT REQUEST IS ACKNOWLEDGED WITH THE REGISTER AT $DA9000. THERE IS NOT A HARDWARE INTERUPT ACK, SO JUST FYI.	
	
	PROCESS (CPUCLK) BEGIN
		IF (RISING_EDGE (CPUCLK)) THEN
		
			IF (RnW = '1' AND nAS = '0' AND nIDEDIS = '1') THEN
			
				CASE A(23 DOWNTO 12) IS
					WHEN x"DE1" => DATAOUT <= x"DF"; --GAYLE_ID is at $DE1000. Return $DF (11011111).
					WHEN x"DAA" => DATAOUT <= x"80"; --INTENA (enable ide interupts) AT $DAA000, Return $80 (10000000).
					WHEN x"DA8" => DATAOUT <= INTRQ & "0000001"; --IDE Device Interrupt Request on data bit 7 at $DA8000.
					WHEN OTHERS => DATAOUT <= (OTHERS => 'Z');
				END CASE;
				
			END IF;
			
		END IF;
	END PROCESS;
	
	--ARE WE IN THE ASSIGNED ADDRESS SPACE FOR THE IDE CONTROLLER?
	--GAYLE IDE ADDRESS SPACE IS $0DA0000 - $0DA3FFF. THE ADDRESS SPACE IS HARD CODED IN GAYLE.
	--SPACE $0DA4000 - $0DA4FFF IS IDE RESERVED. AFAIK IT WAS NEVER IMPLEMENTED.
	--WE CONSIDER BGACK BECAUSE WE DON'T WANT TO RESPOND TO DMA GENERATED ADDRESSES.
	--$DA0 = 110110100000, $da3 = 110110100011
	--IDE_SPACE <= '1' WHEN (A(23 DOWNTO 12) >= x"DA0" AND A(23 DOWNTO 12) <= x"DA3") AND nAS = '0' AND nBGACK = '1' ELSE '0';
	IDE_SPACE <= '1' WHEN A(23 DOWNTO 14) = "1101101000" AND nAS = '0' AND nBGACK = '1' ELSE '0';
	
	--GAYLE SPECS TELL US WHEN THE IDE CHIP SELECT LINES ARE ACTIVE
	
	nCS0 <= '0' 
		WHEN 
			(A(13 DOWNTO 12) = "00" OR A(13 DOWNTO 12) = "10") AND nAS = '0' AND IDE_SPACE = '1' --$0DA0000 TO $0DA0FFF OR $0DA2000 TO $0DA2FFF
		ELSE 
			'1';
			
	nCS1 <= '0' 
		WHEN 
			(A(13 DOWNTO 12) = "01" OR A(13 DOWNTO 12) = "11") AND nAS = '0' AND IDE_SPACE = '1' --$0DA1000 TO $0DA1FFF OR $0DA3000 TO $0DA3FFF
		ELSE 
			'1';
			
	--GAYLE EXPECTS IDE DA2..0 TO BE CONNECTED TO A4..2
	
	DA(0) <= A(2);
	DA(1) <= A(3);
	DA(2) <= A(4);	
	
	--HERE IS THE CONTROLLER INTERFACE
	PROCESS (CPUCLK, nRESET) BEGIN
	
		IF (nRESET = '0') THEN
			--AMIGA HAS RESET, START OVER
			nDIOR <= '1';
			nDIOW <= '1';
			--nDSACK0 <= 'Z';
			nDSACK1 <= 'Z';
			nDTACK <= 'Z';
		
		ELSIF (RISING_EDGE(CPUCLK)) THEN
		
			IF (IDE_SPACE = '1') THEN			
				--WE ARE IN THE IDE ADDRESS SPACE 
				--THE TIMINGS HERE MAY NEED SOME TWEAKING
				
				 IF (nAS = '0') THEN 
					--ADDRESS STROBE IS ASSERTED
				
					IF (RnW = '1') THEN
						--THIS IS A READ
						nDIOR <= '0';
						nDIOW <= '1';
					ELSE
						--THIS IS A WRITE
						--THE GAYLE TIMINGS SAY WRITE SHOULD WAIT ONE CLOCK AFTER LDS/UDS, SO THAT MAY NEED TO BE INCLUDED.
						nDIOR <= '1';
						nDIOW <= '0';
					END IF;
						
					IF (IORDY = '1') THEN
						--IORDY IS ACTIVE HIGH BUT IS CALLED "_WAIT" IN THE GAYLE SPECS. 
						--WHEN HIGH, THE IDE DEVICE IS READY TO TRANSMIT OR RECEIVE DATA. 						
						--SIGNAL 16 BIT PORT TO 68030 OR DTACK WHEN WE ARE IN 68K MODE.
						IF (MODE68K = '0') THEN
							--nDSACK0 <= '1';
							nDSACK1 <= '0';
						ELSE
							nDTACK <= '0';
						END IF;
						
					END IF;
					
				ELSE
				
					--ADDRESS STROBE NOT ASSERTED
					IF (MODE68K = '0') THEN
						--nDSACK0 <= '1';
						nDSACK1 <= '1';
					ELSE
						nDTACK <= '1';
					END IF;
					
				END IF;	
			
			ELSE
			
				--SET IN A "NOP" STATE
				nDIOR <= '1';
				nDIOW <= '1';
				
				--HI Z DSACK/DTACK SO WE DON'T INTERFERE WITH OTHER STUFF ON THE BUS
				IF (MODE68K = '0') THEN
					--nDSACK0 <= 'Z';
					nDSACK1 <= 'Z';
				ELSE
					nDTACK <= 'Z';
				END IF;
					
			END IF;
		
		END IF;
	
	END PROCESS;

	------------------------------
	-- ZORRO 3 MEMORY CONTROLER --
	------------------------------
	
	--ARE WE IN THE Z3 ADDRESS SPACE?
	--WE CONSIDER BGACK BECAUSE WE DON'T WANT TO RESPOND TO DMA GENERATED ADDRESSES, ALTHOUGH THAT SHOULD NEVER HAPPEN HERE BECAUSE
	--24 BIT DMA CANNOT ACCESS THE ZORRO 3 MEMORY SPACE.
	--EXTSEL IS A SIGNAL THAT PREVENTS 68K STATE MACHINE ACTIVITIES IN U600. THIS SHOULD NOT CONSIDER ADDRESS STROBE.
	EXTSEL <= '1' WHEN 
			A(31 DOWNTO 27) = Z3RAM_BASE_ADDR AND nBGACK = '1' AND Z3RAM_CONFIGED = '1' AND FC(2 DOWNTO 0) /= "111" 
		ELSE 
			'0';
	
	--ARE WE ACCESSING THE Z3 MEMORY?
	MEMORY_SPACE <= '1' 
		WHEN 
			EXTSEL = '1' AND nAS = '0'
		ELSE 
			'0';

	--DETERMINE WHAT SPACE IN THE MEMORY WE ARE ACCESSING
	--THIS DETERMINES WHICH PAIR OF SDRAMS WE ARE ACCESSING
	LOW_MEMORY_SPACE <= '1' WHEN A(26) = '0' AND MEMORY_SPACE = '1' ELSE '0';
	HIGH_MEMORY_SPACE <= '1' WHEN A(26) = '1' AND MEMORY_SPACE = '1' ELSE '0';
	
--FOR FUTURE CONSIDERATION...ALLOWING MULTIPLE RAM CONFIGURATIONS UP TO 256MB
--256MB IS THE GREATEST CAPACITY IN THE TSOP 2 PACKAGE. THIS REQUIRES THE ADDITION OF 3 JUMPERS w/PULLUPS TO CONFIGURE.
--So, jumper placed = 0 (GND), no jumper = 1

--RAMSIZE = vector (0..2) (JM0..1..2)
--
--case ramsize
--
--	when "011" then if A(24) = '0' then lowpage else highpage --32MB
--	when "010" then if A(25) = '0' then lowpage else highpage --64MB
--	when "001" then if A(26) = '0' then lowpage else highpage --128MB
--	when "000" then if A(27) = '0' then lowpage else highpage --256MB
--	
--	when others ALWAYS lowpage
--	
--end case
--
--to support 256mb, need to connect through A26 to SDRAM and possibly alter autoconfig
	
	--SET THE DYNAMIC BUS SIZING
	--THIS IS SILLY. COMBINE THESE INTO A SINGLE SET OF OUTPUTS FOR NEXT REVISION.
	nEM0UUBE <= nUUBE;
	nEM0UMBE <= nUMBE;
	nEM0LMBE <= nLMBE;
	nEM0LLBE <= nLLBE;
	
	nEM1UUBE <= nUUBE;
	nEM1UMBE <= nUMBE;
	nEM1LMBE <= nLMBE;
	nEM1LLBE <= nLLBE;
	
	--------------------------------------
	-- SDRAM FALLING CLOCK EDGE ACTIONS --
	--------------------------------------
	
	--ALL THE NECESSARY RAM TIMINGS WITH PAL EQUATIONS ARE IN THE 68030 MANUAL, SECTIONS 7 AND 12
	
	PROCESS ( CPUCLK ) BEGIN
		
		IF ( FALLING_EDGE (CPUCLK) ) THEN

			IF (MEMORY_SPACE = '1') THEN		

				--ENABLE THE VARIOUS BYTES ON THE SDRAM DEPENDING ON WHAT THE ACCESSING DEVICE IS ASKING FOR.
				--DISCUSSION OF PORT SIZE AND BYTE ACTIVATION IS ALL IN SECTION 12 OF THE 68030 USER MANUAL.
				
				--UPPER UPPER BYTE ENABLE (D31..24)
				IF 
				   (( RnW = '1' ) OR
					(A(1 downto 0) = "00" AND nDS = '0'))
				THEN			
					nUUBE <= '0'; 
				ELSE 
					nUUBE <= '1';
				END IF;

				--UPPER MIDDLE BYTE (D23..16)
				IF 
					(( RnW = '1' ) OR
					(A(1 downto 0) = "01" AND nDS = '0') OR
					(A(1) = '0' AND SIZ(0) = '0'  AND nDS = '0') OR
					(A(1) = '0' AND SIZ(1) = '1'  AND nDS = '0')) 
				THEN
					nUMBE <= '0';
				ELSE
					nUMBE <= '1';
				END IF;

				--LOWER MIDDLE BYTE (D15..8)
				IF 
				   (( RnW = '1' ) OR
					(A(1 downto 0) = "10" AND nDS = '0') OR
					(A(1) = '0' AND SIZ(0) = '0' AND SIZ(1) = '0'  AND nDS = '0') OR
					(A(1) = '0' AND SIZ(0) = '1' AND SIZ(1) = '1'  AND nDS = '0') OR
					(A(0) = '1' AND A(1) = '0' AND SIZ(0) = '0'  AND nDS = '0'))
				THEN
					nLMBE <= '0';
				ELSE
					nLMBE <= '1';
				END IF;

				--LOWER LOWER BYTE (D7..0)
				IF 
				   (( RnW = '1' ) OR
					(A(1 downto 0) = "11" AND nDS = '0' ) OR
					(A(0) = '1' AND SIZ(0) = '1' AND SIZ(1) = '1' AND nDS = '0') OR
					(SIZ(0) = '0' AND SIZ(1) = '0' AND nDS = '0') OR
					(A(1) = '1' AND SIZ(1) ='1' AND nDS = '0'))
				THEN
					nLLBE <= '0';
				ELSE
					nLLBE <= '1';
				END IF;	

			ELSE 
				--DEACTIVATE ALL THE RAM BYTE MASKS

				nUUBE <= '1';
				nUMBE <= '1';
				nLMBE <= '1';
				nLLBE <= '1';

			END IF;	
		END IF;
	END PROCESS;
	
	
	-------------------------------------
	-- SDRAM RISING CLOCK EDGE ACTIONS --
	-------------------------------------
	
	PROCESS ( CPUCLK, nGRESET ) BEGIN
	
		IF (nGRESET = '0') THEN 
				--THE AMIGA HAS BEEN RESET
				CURRENT_STATE <= POWERUP;
				
				nCAS0 <= '1';
				nRAS0 <= '1';
				nEM0WE <= '1';
				nEM0CS <= '1';
				EM0CLKE <= '0';
				
				nCAS1 <= '1';
				nRAS1 <= '1';
				nEM1WE <= '1';
				nEM1CS <= '1';
				EM1CLKE <= '0';
				
				COUNT <= 0;
				SDRAM_START_REFRESH_COUNT <= '0';
				nSTERM <= 'Z';
				
		ELSIF ( RISING_EDGE (CPUCLK) ) THEN
			
			--SDRAM is pretty fast. Most operations will complete in less than one 25MHz clock cycle. Only AUTOREFRESH and 
			--successive BANK ACTIVE commands take more than one clock cycle. Both are 60ns.
			
			--NEED TO IMPLEMENT BURST WITH BERR!!!!!!!!!
			
			--REFRESH
			IF (REFRESH_COUNTER >= REFRESH_COUNTER_DEFAULT AND CURRENT_STATE /= DATA_STATE) THEN
				--TIME TO REFRESH THE SDRAM
				IF (MEMORY_SPACE = '0') THEN
					--IF THIS IS NOT A MEMORY CYCLE, PROCEED DIRECTLY TO REFRESH
					--IF WE ARE IN THE MIDDLE OF MEMORY ACCESS, WE NEED TO WAIT UNTIL THAT IS OVER
					CURRENT_STATE <= AUTO_REFRESH;
				END IF;
			ELSE
				--INCREMENT THE REFRESH COUNTER
				REFRESH_COUNTER <= REFRESH_COUNTER + 1;
			END IF;
		
			--PROCEED WITH SDRAM STATE MACHINE
			--THE FIRST STATES ARE TO INITIALIZE THE SDRAM, WHICH WE ALWAYS DO
			--THE LATER STATES ARE TO UTILIZE THE SDRAM, WHICH ONLY HAPPENS IF MEMORY_SPACE = 1
			--THIS MEANS THE ADDRESS STROBE IS ASSERTED, WE ARE IN THE ZORRO 3 ADDRESS SPACE, AND THE RAM IS AUTOCONFIGured
			CASE CURRENT_STATE IS
			
				WHEN POWERUP =>
					--First power up or warm reset
					--200 microsecond is needed to stabilize. We are going to rely on the 
					--the system reset timer to give us the needed time, although it might be inadequate.
					
					nCAS0 <= '1';
					nRAS0 <= '1';
					nEM0WE <= '1';
					nEM0CS <= '1';
					EM0CLKE <= '0';
					
					nCAS1 <= '1';
					nRAS1 <= '1';
					nEM1WE <= '1';
					nEM1CS <= '1';
					EM1CLKE <= '0';
					
					CURRENT_STATE <= POWERUP_PRECHARGE;
					
				WHEN POWERUP_PRECHARGE =>
					--ALL BANKS TO BE PRECHARGED
					EMA <= (OTHERS => '0');
					EMA(10) <= '1'; --PRECHARGE ALL	
					
					nCAS0 <= '1';
					nRAS0 <= '0';
					nEM0WE <= '0';
					nEM0CS <= '0';
					EM0CLKE <= '1';
					
					nCAS1 <= '1';
					nRAS1 <= '0';
					nEM1WE <= '0';
					nEM1CS <= '0';
					EM1CLKE <= '1';
					
					CURRENT_STATE <= MODE_REGISTER;
				
				WHEN MODE_REGISTER =>
					--TWO CLOCK CYCLES ARE NEEDED FOR THE REGISTER TO, WELL, REGISTER
					EMA <= "0001000100000"; --PROGRAM THE SDRAM...NO READ OR WRITE BURST, CAS LATENCY=2,
					
					nCAS0 <= '0';
					nRAS0 <= '0';
					nEM0WE <= '0';
					nEM0CS <= '0';
					
					nCAS1 <= '0';
					nRAS1 <= '0';
					nEM1WE <= '0';
					nEM1CS <= '0';
					
					IF (COUNT = 1) THEN
						--NOW NEED TO REFRESH TWICE
						CURRENT_STATE <= AUTO_REFRESH;
					END IF;
					
					COUNT <= COUNT + 1;
					
				WHEN AUTO_REFRESH =>
					--REFRESH the SDRAM
					--MUST BE FOLLOWED BY NOPs UNTIL REFRESH COMPLETE
					--Refresh time is 60ns. Each 25MHz clock period is 40ns.
					--If we wait two clock cycles, this will allow time for refresh.
					
					nCAS0 <= '0';
					nRAS0 <= '0';
					nEM0WE <= '1';
					nEM0CS <= '0';
					
					nCAS1 <= '0';
					nRAS1 <= '0';
					nEM1WE <= '1';
					nEM1CS <= '0';					
					
					COUNT <= 0;
					
					CURRENT_STATE <= AUTO_REFRESH_CYCLE;				
					
				WHEN AUTO_REFRESH_CYCLE =>
					--NOPs WHILE THE SDRAM IS REFRESHING
					
					nCAS0 <= '1';
					nRAS0 <= '1';
					nEM0WE <= '1';
					nEM0CS <= '0';
					
					nCAS1 <= '1';
					nRAS1 <= '1';
					nEM1WE <= '1';
					nEM1CS <= '0';	
					
					--IF (COUNT = 1) THEN --TWO CLOCK CYCLES HAVE PASSED. WE CAN PROCEED.
						--I THINK THIS IS AN EXTRA CLOCK CYCLE BECAUSE THE PREVIOUS CLOCK CYCLE SHOULD BE INCLUDED IN THE COUNT
						--DO WE NEED TO REFRESH AGAIN (BECAUSE WE'RE STILL IN STARTUP CONDITIONS)?
						IF (SDRAM_START_REFRESH_COUNT = '0') THEN							
							CURRENT_STATE <= AUTO_REFRESH;
							SDRAM_START_REFRESH_COUNT <= '1';
						ELSE
							--DESELECT ALL SDRAMs
							nEM0CS <= '1';
							nEM1CS <= '1';	
							
							--WE SHOULD BE READY TO GO!
							CURRENT_STATE <= RUN_STATE;
							REFRESH_COUNTER <= 0;
						END IF;
					--END IF;		

					COUNT <= COUNT + 1;						
				
				WHEN RUN_STATE =>
					--CLOCK EDGE 0
					
					IF (MEMORY_SPACE = '1') THEN 
						--WE ARE IN THE Z3 MEMORY SPACE WITH THE ADDRESS STROBE ASSERTED.
						--SEND THE BANK ACTIVATE COMMAND W/RAS
						
						--SELECT THE CORRECT SET OF SDRAMs BASED ON ADDRESS
						IF (LOW_MEMORY_SPACE = '1') THEN nEM0CS <= '0'; ELSE nEM0CS <= '1'; END IF;
						IF (HIGH_MEMORY_SPACE = '1') THEN nEM1CS <= '0'; ELSE nEM1CS <= '1'; END IF;
						
						EMA(12 downto 0) <= A(14 downto 2);
						BANK0 <= A(15);
						BANK1 <= A(16);
						
						--HERE, I'M SENDING THE COMMANDS TO ALL SDRAMs, BUT ONLY THE SELECTED PAIR SHOULD RESPOND
						nCAS0 <= '1';
						nRAS0 <= '0';
						nEM0WE <= '1';
						
						nCAS1 <= '1';
						nRAS1 <= '0';
						nEM1WE <= '1';
						
						nSTERM <= '1'; --WE ARE USING THE BUS RIGHT NOW, SO NEGATE STERM IN PREPARTATION FOR USE
						
						CURRENT_STATE <= CAS_STATE;
						COUNT <= 0;
					END IF;
					
				WHEN CAS_STATE =>
					--CLOCK EDGE 1
					--READ OR WRITE WITH AUTOPRECHARGE
					
					EMA(8 downto 0) <= A(25 downto 17);
					EMA(9) <= '0';
					EMA(10) <= '1'; --AUTO PRECHARGE
					
					nCAS0 <= '0';
					nRAS0 <= '1';
					nEM0WE <= RnW;
					
					nCAS1 <= '0';
					nRAS1 <= '1';
					nEM1WE <= RnW;

					--IF THIS IS A WRITE ACTION, WE CAN IMMEDIATELY PROCEED TO THE ACTION
					--IF THIS IS A READ ACTION, THE CAS LATENCY IS 2 CLOCK CYCLES, SO WE NEED TO WAIT ONE MORE CLOCK BEFORE READING
					--DATA STROBE IS NOT REALLY NEEDED WITH WRITE EVENTS

					IF ((RnW = '0') OR (RnW = '1' AND COUNT >= 1 AND nDS = '0')) THEN
					
						nSTERM <= '0';
						
						CURRENT_STATE <= DATA_STATE;
					
					END IF;						
					
					COUNT <= COUNT + 1;
					
				WHEN DATA_STATE =>
					--RISING CLOCK EDGE 2
					--THIS IS THE CLOCK EDGE WE EXPECT THE DATA TO BE WRITTEN TO OR READ FROM THE SDRAM
					--WE NEED TO WAIT 30ns BEFORE ISSUING ANOTHER BANK ACTIVATE COMMAND. NO PROBLEM, SINCE ONE CLOCK CYCLE IS 40ns.
					
					IF (MEMORY_SPACE = '0') THEN --THE ADDRESS STROBE HAS NEGATED INDICATING THE END OF THE MEMORY ACCESS
						
						--TRISTATE SO WE DON'T INTERFERE WITH OTHER DEVICES ON THE BUS
						nSTERM <= 'Z';
						
						CURRENT_STATE <= RUN_STATE;
						
						--SET NOP
						nCAS0 <= '1';
						nRAS0 <= '1';
						nEM0WE <= '1';
						nEM0CS <= '1';
						
						nCAS1 <= '1';
						nRAS1 <= '1';
						nEM1WE <= '1';
						nEM1CS <= '1';
						
					END IF;					
				
			END CASE;
				
		END IF;
	END PROCESS;

end Behavioral;

